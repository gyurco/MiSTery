// vidclkcntrl.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module vidclkcntrl (
		input  wire  inclk1x,   //  altclkctrl_input.inclk1x
		input  wire  inclk0x,   //                  .inclk0x
		input  wire  clkselect, //                  .clkselect
		output wire  outclk     // altclkctrl_output.outclk
	);

	vidclkcntrl_altclkctrl_0 altclkctrl_0 (
		.inclk1x   (inclk1x),   //  altclkctrl_input.inclk1x
		.inclk0x   (inclk0x),   //                  .inclk0x
		.clkselect (clkselect), //                  .clkselect
		.outclk    (outclk)     // altclkctrl_output.outclk
	);

endmodule
