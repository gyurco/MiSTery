//
// audio.v
// 
// Atari audio subsystem implementation for the MiST board
// http://code.google.com/p/mist-board/
// 
// Copyright (c) 2015 Till Harbaum <till@harbaum.org> 
// 
// This source file is free software: you can redistribute it and/or modify 
// it under the terms of the GNU General Public License as published 
// by the Free Software Foundation, either version 3 of the License, or 
// (at your option) any later version. 
// 
// This source file is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the 
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License 
// along with this program.  If not, see <http://www.gnu.org/licenses/>. 

module audio (
	// system interface
	input  	reset,
	input 	clk,      // 32 MHz
	input   clk_8_en,
	input   clk_2_en,
	input [1:0] bus_cycle,   // bus-cycle for sync
	

	// cpu interface
	input [15:0] din,
	input [15:0] addr,
	output [15:0] dout,
	input uds,
	input lds,
	input rw,
	input psg_sel,
	input ste_dma_snd_sel,

	// ste dma interface
	input			hde1,     // to synchronize with video
	output            dma_read,
	output [22:0]     dma_addr,
	input [63:0]      dma_data,
	
	input psg_stereo,
	
	// psg has gpios
	output floppy_side,
	output [1:0] floppy_sel,
	// extra joystick map to parallel port
	input [5:0] joy0,
	input [5:0] joy1,
	
	output [7:0] parallel_data_out,
	input parallel_strobe_out,
	output parallel_data_out_available,
	
	output 				xsint,
	output 				xsint_d,
	
	output audio_r,
	output audio_l
);
	
wire [7:0] port_a_out;
wire [7:0] port_b_out;
assign floppy_side = port_a_out[0];
assign floppy_sel = port_a_out[2:1];

wire [9:0] ym_audio_out_l, ym_audio_out_r;
wire [7:0] ym_a_out, ym_b_out, ym_c_out;

assign ym_audio_out_l = psg_stereo ? ym_a_out + ym_b_out : ym_a_out + ym_b_out + ym_c_out;
assign ym_audio_out_r = psg_stereo ? ym_c_out + ym_b_out : ym_a_out + ym_b_out + ym_c_out;

// extra joysticks are wired to the printer port
// using the "gauntlet2 interface", fire of 
// joystick 0 is connected to the mfp I0 (busy)
wire [7:0] port_b_in = { ~joy0[0], ~joy0[1], ~joy0[2], ~joy0[3], 
								 ~joy1[0], ~joy1[1], ~joy1[2], ~joy1[3]}; 
wire [7:0] port_a_in = { 2'b11, ~joy1[4], 5'b11111 }; 

assign dout = psg_sel?{psg_dout,8'hff}:ste_dma_snd_sel?ste_dma_snd_data_out:16'h0000;
wire [15:0] ste_dma_snd_data_out;
wire [7:0] psg_dout;

ym2149 ym2149 (
	.CLK         ( clk                ),
	.CE          ( clk_2_en           ),
	.RESET       ( reset              ),
	.DI          ( din[15:8]          ),
	.DO          ( psg_dout           ),
	.CHANNEL_A   ( ym_a_out           ),
	.CHANNEL_B   ( ym_b_out           ),
	.CHANNEL_C   ( ym_c_out           ),
	.BDIR        ( psg_sel & ~rw      ),
	.BC          ( psg_sel & ~addr[1] ),
	.MODE        ( 0                  ),
	.SEL         ( 0                  ),
	.IOA_in      ( port_a_in          ),
	.IOA_out     ( port_a_out         ),
	.IOB_in      ( port_b_in          ),
	.IOB_out     ( port_b_out         )
);
wire parallel_fifo_full;

// ------ fifo to store printer data coming from psg ---------
io_fifo #(.DEPTH(4)) parallel_out_fifo (
	.reset 				(reset),		

	.in_clk  			(clk),
	.in 				(port_b_out),
	.in_strobe 			(port_a_out[5]),
	.in_enable		 	(1'b0),

	.out_clk  			(clk),
	.out 				(parallel_data_out),
	.out_strobe 		(parallel_strobe_out),
	.out_enable		 	(1'b0),

	.full					(parallel_fifo_full),
	.data_available 	(parallel_data_out_available)
);

wire [7:0] ste_audio_out_r;
wire [7:0] ste_audio_out_l;

ste_dma_snd ste_dma_snd (
	// cpu interface
	.clk        (clk             ),
	.clk_8_en   (clk_8_en        ),
	.reset      (reset           ),
	.din        (din             ),
	.sel        (ste_dma_snd_sel ),
	.addr       (addr[5:1]       ),
	.uds        (uds             ),
	.lds        (lds             ),
	.rw         (rw              ),
	.dout       (ste_dma_snd_data_out),

	// memory interface
	.clk_2_en   (clk_2_en        ),
	.bus_cycle 	(bus_cycle       ),
	.hde1       (hde1            ),
	.saddr      (dma_addr        ),
	.read       (dma_read        ),
	.data       (dma_data        ),

	.audio_l    (ste_audio_out_l ),
	.audio_r    (ste_audio_out_r ),

	.xsint     	( xsint ),
	.xsint_d   	( xsint_d )   // 4 usec delayed
);

// audio output processing

// YM and STE audio channels are expanded to 14 bits and added resulting in 15 bits 
// for the sigmadelta dac take from the minimig

// This should later be handled by the lmc1992

wire [9:0] ym_audio_out_l_signed = ym_audio_out_l - 10'h200;
wire [9:0] ym_audio_out_r_signed = ym_audio_out_r - 10'h200;
wire [7:0] ste_audio_out_l_signed = ste_audio_out_l - 8'h80;
wire [7:0] ste_audio_out_r_signed = ste_audio_out_r - 8'h80;

wire [14:0] audio_mix_l = 
	{ ym_audio_out_l_signed[9], ym_audio_out_l_signed, ym_audio_out_l_signed[9:6]} + 
	{ ste_audio_out_l_signed[7], ste_audio_out_l_signed, ste_audio_out_l_signed[7:2] };
wire [14:0] audio_mix_r = 
	{ ym_audio_out_r_signed[9], ym_audio_out_r_signed, ym_audio_out_r_signed[9:6]} + 
	{ ste_audio_out_r_signed[7], ste_audio_out_r_signed, ste_audio_out_r_signed[7:2] };

sigma_delta_dac sigma_delta_dac (
	.clk      ( clk         ),	// bus clock
	.ldatasum ( audio_mix_l ),	// left channel data
	.rdatasum ( audio_mix_r ),	// right channel data
	.left   	 ( audio_l     ),	// left bitstream output
	.right	 ( audio_r     )	// right bitsteam output
);

endmodule
